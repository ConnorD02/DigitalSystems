module mulTB;

logic